`timescale 1ns / 1ps
/*
fwdcombine.v

The complement to snoopsplit 
*/


module fwdcombine(

    );
endmodule

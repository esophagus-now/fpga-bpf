`timescale 1ns / 1ps
/*
snoop_arbiter_3.v

The "3" in the name was chosen because it has three inputs, but I probably
should have called it snoop_arbiter_2.v, since the "any_in" input is more
of like a "carry in". Oh well

A primitive used inside parallel_packetfilts.v. Essentially, this ends up
deciding which of the packet filters will receive data from the snooper,
depending on which ones are ready.

This module was carefully written in order to have the minimum combinational
delay. I went back and forth between editing the Verilog and looking at the 
synthesized circuit generated by Vivado.
*/


module snoop_arbiter_3(
	input wire any_in,
	input wire mem_ready_left,
	input wire mem_ready_right,
	output wire en_left,
	output wire en_right,
	output wire any_out
);

assign en_left = !any_in && mem_ready_left;
assign en_right = !any_in && !mem_ready_left && mem_ready_right;
assign any_out = any_in || mem_ready_left || mem_ready_right;

endmodule

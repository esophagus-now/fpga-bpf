`timescale 1ns / 1ps
/*
snoop_arbiter_5.v

The "5" in the name was chosen because it has five inputs, but I probably
should have called it snoop_arbiter_4.v, since the "any_in" input is more
of like a "carry in". Oh well

A primitive used inside parallel_packetfilts.v. Essentially, this ends up
deciding which of the packet filters will receive data from the snooper,
depending on which ones are ready.

This module was carefully written in order to have the minimum combinational
delay. I went back and forth between editing the Verilog and looking at the 
synthesized circuit generated by Vivado.
*/

//Yes I'm the arbiter my word is law-aw-aw...
module arbiter_4 (
	input wire any_in,
	input wire mem_ready_A,
	input wire mem_ready_B,
	input wire mem_ready_C,
	input wire mem_ready_D,
	output wire en_A,
	output wire en_B,
	output wire en_C,
	output wire en_D,
	output wire any_out
);

assign en_A = !any_in && mem_ready_A;
assign en_B = !any_in && !mem_ready_A && mem_ready_B;
assign en_C = !any_in && !mem_ready_A && !mem_ready_B && mem_ready_C;
assign en_D = !any_in && !mem_ready_A && !mem_ready_B && !mem_ready_C && mem_ready_D;
assign any_out = any_in || mem_ready_A || mem_ready_B || mem_ready_C || mem_ready_D;

endmodule
